module and_gate(in1, in2, out);
input in1, in2;
output out;
and(out, in1, in2);
endmodule

