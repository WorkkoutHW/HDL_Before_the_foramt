module prog_mem(addr, dout);

	input	[7:0]	addr;
	output	[15:0]	dout;

	reg 	[15:0]	rom[0:255];

	assign 	dout = rom[addr];

initial
	begin
		rom[8'h00] = 16'b1100_0001_0010_0000;  	//LDI $value R0
		rom[8'h01] = 16'b1100_0011_0100_0001;  	//LDI $value R1
		rom[8'h02] = 16'b1100_0101_0110_0010;  	//LDI $value R2
		rom[8'h03] = 16'b1100_0111_1000_1100;  	//LDI $value R12
		rom[8'h04] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h05] = 16'b0001_0000_0001_0100;  	//ADD R0 R1 R4
		rom[8'h06] = 16'b0010_0000_0001_0101; 	//SUB R0 R1 R5 
		rom[8'h07] = 16'b0011_0000_xxxx_0000; 	//DEC R0    R0 
		rom[8'h08] = 16'b0100_0000_0001_0010;  	//AND R0 R1 R2
		rom[8'h09] = 16'b0101_0000_0001_0010;  	//IOR R0 R1 R2
		rom[8'h0a] = 16'b0110_0000_0001_0010;  	//XOR R0 R1 R2
		rom[8'h0b] = 16'b0111_0000_xxxx_0010;  	//INV R0    R2
		rom[8'h0c] = 16'b1000_0000_xxxx_0000;  	//SHR R0    R0
		rom[8'h0d] = 16'b1001_0001_xxxx_0001;   //SHL R1    R1
		rom[8'h0e] = 16'b1010_0100_xxxx_0010;  	//MOV R4    R2
		rom[8'h0f] = 16'b1100_0001_0011_1111;  	//JUI $value	(LDI $value R15)
		rom[8'h10] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h11] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h12] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h13] = 16'b1100_1111_1111_0001;  	//LDI $value R1
		rom[8'h14] = 16'b1100_0000_0001_0010;  	//LDI $value R2
		rom[8'h15] = 16'b0001_0001_0010_0010; 	//ADD R1 R2 R2 
		rom[8'h16] = 16'b1110_xxxx_xxxx_1000;  	//JES 
		rom[8'h17] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h18] = 16'b1110_xxxx_xxxx_0100;  	//JFS
		rom[8'h19] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h1a] = 16'b1110_0000_0000_0001;  	//JEQ R0 R0
		rom[8'h1b] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0
		rom[8'h1c] = 16'b1111_xxxx_xxxx_0010; 	//CLE 
		rom[8'h1d] = 16'b1111_xxxx_0000_0100;  	//VMW    R0		
		rom[8'h1e] = 16'b1111_xxxx_0001_1000; 	//DMW 	 R1
		rom[8'h1f] = 16'b1101_xxxx_xxxx_0110;  	//DMR	    R6
		rom[8'h20] = 16'b1010_1111_xxxx_1111;  	//JUD R2  	(MOV R2    R15)
		rom[8'h21] = 16'b0000_0000_xxxx_0000;  	//INC R0    R0  	
		rom[8'h22] = 16'bxxxx_xxxx_xxxx_xxxx;  	
		rom[8'h23] = 16'bxxxx_xxxx_xxxx_xxxx;  	
		rom[8'h24] = 16'bxxxx_xxxx_xxxx_xxxx;  	
		rom[8'h25] = 16'bxxxx_xxxx_xxxx_xxxx;  	
		rom[8'h26] = 16'bxxxx_xxxx_xxxx_xxxx;	
		rom[8'h27] = 16'b0000_0000_0000_0000;  	
		rom[8'h28] = 16'b1111_0000_0000_0010;  	
		rom[8'h29] = 16'b0000_0000_0000_0000;  	
		rom[8'h2a] = 16'b1111_0000_0000_0001;  	
		rom[8'h2b] = 16'b0000_0000_0000_0000;  	
		rom[8'h2c] = 16'b1110_0100_0000_0000; 	 
		rom[8'h2d] = 16'b1110_0010_0000_0000;  			
		rom[8'h2e] = 16'b1110_0001_0001_0000; 	
		rom[8'h2f] = 16'b1101_0000_0000_0110;  	
		rom[8'h30] = 16'b1100_0001_0010_0000;  	
		rom[8'h31] = 16'b1100_0011_0100_0001;  	
		rom[8'h32] = 16'b1100_0101_0110_0010;  	
		rom[8'h33] = 16'b1100_0111_1000_1100;  	
		rom[8'h34] = 16'b0000_0000_0000_0000;  	
		rom[8'h35] = 16'b0001_0000_0001_0100;  	
		rom[8'h36] = 16'b0010_0000_0001_0101; 	 
		rom[8'h37] = 16'b0011_0000_0000_0000; 	 
		rom[8'h38] = 16'b0100_0000_0001_0010;  	
		rom[8'h39] = 16'b0101_0000_0001_0010;  	
		rom[8'h3a] = 16'b0110_0000_0001_0010;  	
		rom[8'h3b] = 16'b0111_0000_0000_0010;  	
		rom[8'h3c] = 16'b1000_0000_0000_0000;  	
		rom[8'h3d] = 16'b1001_0001_0000_0001;   
		rom[8'h3e] = 16'b1010_0100_0000_0010;  	
		rom[8'h3f] = 16'b1100_0001_0011_1111;  		
		rom[8'h40] = 16'b0000_0000_0000_0000;  	
		rom[8'h41] = 16'b0000_0000_0000_0000;  	
		rom[8'h42] = 16'b0000_0000_0000_0000;  	
		rom[8'h43] = 16'b1100_1111_1111_0001;  	
		rom[8'h44] = 16'b1100_0000_0001_0010;  	
		rom[8'h45] = 16'b0001_0001_0010_0010; 	 
		rom[8'h46] = 16'b1111_0000_0000_0100;  	
		rom[8'h47] = 16'b0000_0000_0000_0000;  	
		rom[8'h48] = 16'b1111_0000_0000_0010;  	
		rom[8'h49] = 16'b0000_0000_0000_0000;  	
		rom[8'h4a] = 16'b1111_0000_0000_0001;  	
		rom[8'h4b] = 16'b0000_0000_0000_0000;  	
		rom[8'h4c] = 16'b1110_0100_0000_0000; 	 
		rom[8'h4d] = 16'b1110_0010_0000_0000;  		
		rom[8'h4e] = 16'b1110_0001_0001_0000; 	
		rom[8'h4f] = 16'b1101_0000_0000_0110;  	
		rom[8'h50] = 16'b1100_0001_0010_0000;  	
		rom[8'h51] = 16'b1100_0011_0100_0001;  	
		rom[8'h52] = 16'b1100_0101_0110_0010;  	
		rom[8'h53] = 16'b1100_0111_1000_1100;  	
		rom[8'h54] = 16'b0000_0000_0000_0000;  	
		rom[8'h55] = 16'b0001_0000_0001_0100;  	
		rom[8'h56] = 16'b0010_0000_0001_0101; 	
		rom[8'h57] = 16'b0011_0000_0000_0000; 	
		rom[8'h58] = 16'b0100_0000_0001_0010;  	
		rom[8'h59] = 16'b0101_0000_0001_0010;  	
		rom[8'h5a] = 16'b0110_0000_0001_0010;  	
		rom[8'h5b] = 16'b0111_0000_0000_0010;  	
		rom[8'h5c] = 16'b1000_0000_0000_0000;  	
		rom[8'h5d] = 16'b1001_0001_0000_0001;   
		rom[8'h5e] = 16'b1010_0100_0000_0010;  	
		rom[8'h5f] = 16'b1100_0001_0011_1111;  	
		rom[8'h60] = 16'b0000_0000_0000_0000;  	
		rom[8'h61] = 16'b0000_0000_0000_0000;  	
		rom[8'h62] = 16'b0000_0000_0000_0000;  	
		rom[8'h63] = 16'b1100_1111_1111_0001;  	
		rom[8'h64] = 16'b1100_0000_0001_0010;  	
		rom[8'h65] = 16'b0001_0001_0010_0010; 	
		rom[8'h66] = 16'b1111_0000_0000_0100;  	
		rom[8'h67] = 16'b0000_0000_0000_0000;  	
		rom[8'h68] = 16'b1111_0000_0000_0010;  	
		rom[8'h69] = 16'b0000_0000_0000_0000;  	
		rom[8'h6a] = 16'b1111_0000_0000_0001;  	
		rom[8'h6b] = 16'b0000_0000_0000_0000;  	
		rom[8'h6c] = 16'b1110_0100_0000_0000; 	
		rom[8'h6d] = 16'b1110_0010_0000_0000;  		
		rom[8'h6e] = 16'b1110_0001_0001_0000; 	
		rom[8'h6f] = 16'b1101_0000_0000_0110;  	
		rom[8'h70] = 16'b1100_0001_0010_0000;  	
		rom[8'h71] = 16'b1100_0011_0100_0001;  	
		rom[8'h72] = 16'b1100_0101_0110_0010;  	
		rom[8'h73] = 16'b1100_0111_1000_1100;  	
		rom[8'h74] = 16'b0000_0000_0000_0000;  	
		rom[8'h75] = 16'b0001_0000_0001_0100;  	
		rom[8'h76] = 16'b0010_0000_0001_0101; 	
		rom[8'h77] = 16'b0011_0000_0000_0000; 	
		rom[8'h78] = 16'b0100_0000_0001_0010;  	
		rom[8'h79] = 16'b0101_0000_0001_0010;  	
		rom[8'h7a] = 16'b0110_0000_0001_0010;  	
		rom[8'h7b] = 16'b0111_0000_0000_0010;  	
		rom[8'h7c] = 16'b1000_0000_0000_0000;  	
		rom[8'h7d] = 16'b1001_0001_0000_0001;   
		rom[8'h7e] = 16'b1010_0100_0000_0010;  	
		rom[8'h7f] = 16'b1100_0001_0011_1111;  	
		rom[8'h80] = 16'b1100_0001_0010_0000;  	
		rom[8'h81] = 16'b1100_0011_0100_0001;  	
		rom[8'h82] = 16'b1100_0101_0110_0010;  	
		rom[8'h83] = 16'b1100_0111_1000_1100;  	
		rom[8'h84] = 16'b0000_0000_0000_0000;  	
		rom[8'h85] = 16'b0001_0000_0001_0100;  	
		rom[8'h86] = 16'b0010_0000_0001_0101; 	
		rom[8'h87] = 16'b0011_0000_0000_0000; 	
		rom[8'h88] = 16'b0100_0000_0001_0010;  	
		rom[8'h89] = 16'b0101_0000_0001_0010;  	
		rom[8'h8a] = 16'b0110_0000_0001_0010;  	
		rom[8'h8b] = 16'b0111_0000_0000_0010;  	
		rom[8'h8c] = 16'b1000_0000_0000_0000;  	
		rom[8'h8d] = 16'b1001_0001_0000_0001;   
		rom[8'h8e] = 16'b1010_0100_0000_0010;  	
		rom[8'h8f] = 16'b1100_0001_0011_1111;  	
		rom[8'h90] = 16'b0000_0000_0000_0000;  	
		rom[8'h91] = 16'b0000_0000_0000_0000;  	
		rom[8'h92] = 16'b0000_0000_0000_0000;  	
		rom[8'h93] = 16'b1100_1111_1111_0001;  	
		rom[8'h94] = 16'b1100_0000_0001_0010;  	
		rom[8'h95] = 16'b0001_0001_0010_0010; 	
		rom[8'h96] = 16'b1111_0000_0000_0100;  	
		rom[8'h97] = 16'b0000_0000_0000_0000;  	
		rom[8'h98] = 16'b1111_0000_0000_0010;  	
		rom[8'h99] = 16'b0000_0000_0000_0000;  	
		rom[8'h9a] = 16'b1111_0000_0000_0001;  	
		rom[8'h9b] = 16'b0000_0000_0000_0000;  	
		rom[8'h9c] = 16'b1110_0100_0000_0000; 	
		rom[8'h9d] = 16'b1110_0010_0000_0000;  		
		rom[8'h9e] = 16'b1110_0001_0001_0000; 	
		rom[8'h9f] = 16'b1101_0000_0000_0110;  	
		rom[8'ha0] = 16'b1100_0001_0010_0000;  	
		rom[8'ha1] = 16'b1100_0011_0100_0001;  	
		rom[8'ha2] = 16'b1100_0101_0110_0010;  	
		rom[8'ha3] = 16'b1100_0111_1000_1100;  	
		rom[8'ha4] = 16'b0000_0000_0000_0000;  	
		rom[8'ha5] = 16'b0001_0000_0001_0100;  	
		rom[8'ha6] = 16'b0010_0000_0001_0101; 	 
		rom[8'ha7] = 16'b0011_0000_0000_0000; 	
		rom[8'ha8] = 16'b0100_0000_0001_0010;  	
		rom[8'ha9] = 16'b0101_0000_0001_0010;  	
		rom[8'haa] = 16'b0110_0000_0001_0010;  	
		rom[8'hab] = 16'b0111_0000_0000_0010;  	
		rom[8'hac] = 16'b1000_0000_0000_0000;  	
		rom[8'had] = 16'b1001_0001_0000_0001;   
		rom[8'hae] = 16'b1010_0100_0000_0010;  	
		rom[8'haf] = 16'b1100_0001_0011_1111;  	
		rom[8'hb0] = 16'b0000_0000_0000_0000;  	
		rom[8'hb1] = 16'b0000_0000_0000_0000;  	
		rom[8'hb2] = 16'b0000_0000_0000_0000;  	
		rom[8'hb3] = 16'b1100_1111_1111_0001;  	
		rom[8'hb4] = 16'b1100_0000_0001_0010;  	
		rom[8'hb5] = 16'b0001_0001_0010_0010; 	 
		rom[8'hb6] = 16'b1111_0000_0000_0100;  	 
		rom[8'hb7] = 16'b0000_0000_0000_0000;  	
		rom[8'hb8] = 16'b1111_0000_0000_0010;  	
		rom[8'hb9] = 16'b0000_0000_0000_0000;  	
		rom[8'hba] = 16'b1111_0000_0000_0001;  	
		rom[8'hbb] = 16'b0000_0000_0000_0000;  	
		rom[8'hbc] = 16'b1110_0100_0000_0000; 	
		rom[8'hbd] = 16'b1110_0010_0000_0000;  		
		rom[8'hbe] = 16'b1110_0001_0001_0000; 	
		rom[8'hbf] = 16'b1101_0000_0000_0110;  	
		rom[8'hc0] = 16'b1100_0001_0010_0000;  	
		rom[8'hc1] = 16'b1100_0011_0100_0001;  	
		rom[8'hc2] = 16'b1100_0101_0110_0010;  	
		rom[8'hc3] = 16'b1100_0111_1000_1100;  	
		rom[8'hc4] = 16'b0000_0000_0000_0000;  	
		rom[8'hc5] = 16'b0001_0000_0001_0100;  	
		rom[8'hc6] = 16'b0010_0000_0001_0101; 	
		rom[8'hc7] = 16'b0011_0000_0000_0000; 	 
		rom[8'hc8] = 16'b0100_0000_0001_0010;  	
		rom[8'hc9] = 16'b0101_0000_0001_0010;  	
		rom[8'hca] = 16'b0110_0000_0001_0010;  	
		rom[8'hcb] = 16'b0111_0000_0000_0010;  	
		rom[8'hcc] = 16'b1000_0000_0000_0000;  	
		rom[8'hcd] = 16'b1001_0001_0000_0001;   
		rom[8'hce] = 16'b1010_0100_0000_0010;  	
		rom[8'hcf] = 16'b1100_0001_0011_1111;  	
		rom[8'hd0] = 16'b0000_0000_0000_0000;  	
		rom[8'hd1] = 16'b0000_0000_0000_0000;  	
		rom[8'hd2] = 16'b0000_0000_0000_0000;  	
		rom[8'hd3] = 16'b1100_1111_1111_0001;  	
		rom[8'hd4] = 16'b1100_0000_0001_0010;  	
		rom[8'hd5] = 16'b0001_0001_0010_0010; 	
		rom[8'hd6] = 16'b1111_0000_0000_0100;  	
		rom[8'hd7] = 16'b0000_0000_0000_0000;  	
		rom[8'hd8] = 16'b1111_0000_0000_0010;  	
		rom[8'hd9] = 16'b0000_0000_0000_0000;  	
		rom[8'hda] = 16'b1111_0000_0000_0001;  	
		rom[8'hdb] = 16'b0000_0000_0000_0000;  	
		rom[8'hdc] = 16'b1110_0100_0000_0000; 	
		rom[8'hdd] = 16'b1110_0010_0000_0000;  		
		rom[8'hde] = 16'b1110_0001_0001_0000; 	
		rom[8'hdf] = 16'b1101_0000_0000_0110;  	
		rom[8'he0] = 16'b1100_0001_0010_0000;  	
		rom[8'he1] = 16'b1100_0011_0100_0001;  	
		rom[8'he2] = 16'b1100_0101_0110_0010;  	
		rom[8'he3] = 16'b1100_0111_1000_1100;  	
		rom[8'he4] = 16'b0000_0000_0000_0000;  	
		rom[8'he5] = 16'b0001_0000_0001_0100;  	
		rom[8'he6] = 16'b0010_0000_0001_0101; 	 
		rom[8'he7] = 16'b0011_0000_0000_0000; 	
		rom[8'he8] = 16'b0100_0000_0001_0010;  	
		rom[8'he9] = 16'b0101_0000_0001_0010;  	
		rom[8'hea] = 16'b0110_0000_0001_0010;  	
		rom[8'heb] = 16'b0111_0000_0000_0010;  	
		rom[8'hec] = 16'b1000_0000_0000_0000;  	
		rom[8'hed] = 16'b1001_0001_0000_0001;   
		rom[8'hee] = 16'b1010_0100_0000_0010;  	
		rom[8'hef] = 16'b1100_0001_0011_1111;  	
		rom[8'hf0] = 16'b0000_0000_0000_0000;  	
		rom[8'hf1] = 16'b0000_0000_0000_0000;  	
		rom[8'hf2] = 16'b0000_0000_0000_0000;  	
		rom[8'hf3] = 16'b1100_1111_1111_0001;  	
		rom[8'hf4] = 16'b1100_0000_0001_0010;  	
		rom[8'hf5] = 16'b0001_0001_0010_0010; 	
		rom[8'hf6] = 16'b1111_0000_0000_0100;  	
		rom[8'hf7] = 16'b0000_0000_0000_0000;  	
		rom[8'hf8] = 16'b1111_0000_0000_0010;  	
		rom[8'hf9] = 16'b0000_0000_0000_0000;  	
		rom[8'hfa] = 16'b1111_0000_0000_0001;  	
		rom[8'hfb] = 16'b0000_0000_0000_0000;  	
		rom[8'hfc] = 16'b1110_0100_0000_0000; 	
		rom[8'hfd] = 16'b1110_0010_0000_0000;  		
		rom[8'hfe] = 16'b1110_0001_0001_0000; 	
		rom[8'hff] = 16'b1101_0000_0000_0110;  	
	end
/*
initial
	begin
		$readmemb("./rom.bin",rom);
	end
*/
/*
always@(*)
case(addr)
8'h00: 	dout = 16'b1100_0001_0010_0000; //LDI $value R0
default:dout = 16'bxxxx_xxxx_xxxx_xxxx;
endcase
*/
endmodule
